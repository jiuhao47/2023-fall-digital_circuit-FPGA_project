module divider
(
    input clk,rstn,
    output cnt_20b
);

endmodule